<svg xmlns="http://www.w3.org/2000/svg" width="480" height="120" viewBox="0 0 480 120">
  <!-- Background transparent -->
  <!-- Icon: stylized W in purple with motion swoosh -->
  <g transform="translate(10,10)">
    <defs>
      <linearGradient id="g1" x1="0" x2="1" y1="0" y2="1">
        <stop offset="0" stop-color="#8B5CF6"/>
        <stop offset="1" stop-color="#6D28D9"/>
      </linearGradient>
    </defs>

    <!-- Circle background -->
    <circle cx="50" cy="50" r="40" fill="url(#g1)"/>

    <!-- W mark -->
    <path d="M28 48 L38 24 L48 56 L60 20 L72 48" fill="none" stroke="#FFFFFF" stroke-width="6" stroke-linecap="round" stroke-linejoin="round"/>

    <!-- small swoosh to indicate motion -->
    <path d="M78 74 C96 68, 110 60, 130 56" fill="none" stroke="#1E293B" stroke-width="4" stroke-linecap="round" opacity="0.08"/>

    <!-- Text -->
    <g transform="translate(120,34)">
      <text x="0" y="0" font-family="Inter, Roboto, Arial, sans-serif" font-weight="700" font-size="36" fill="#1E293B">Wizex</text>
      <text x="0" y="36" font-family="Inter, Roboto, Arial, sans-serif" font-weight="600" font-size="18" fill="#374151">Remit</text>
    </g>
  </g>
</svg>
